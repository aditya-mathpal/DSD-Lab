module Q2(g,b);
	input [3:0]g;
	output reg [3:0]b;
